interface comp_int;
  logic [31:0] a, b;
  logic [0:0] eq, lt, gt;
endinterface

class comp_tx;
  rand bit [31:0] a, b;  
  bit [0:0] eq, lt, gt;
endclass
class comp_cfg;
  
  static virtual comp_int vif;
  
  static mailbox gen2bfm = new();
  static mailbox mon2ckr = new();
  static mailbox mon2cov = new();
  
endclass

program comp_tb;
  comp_env env = new();

  initial begin
    env.run(); 
  end
endprogram
